package shared_pkg;
	integer correct_count = 0 ;
	integer error_count = 0 ;
	bit test_finished ;
endpackage : shared_pkg